function logic f (input a);
  return a;
endfunction
