module m #(
  localparam int MyParam = 1
);
endmodule

