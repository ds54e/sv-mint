`default_nettype none

module module_names_lower_snake_good;
endmodule

`default_nettype wire
