module m;
endmodule

