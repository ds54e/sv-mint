`default_nettype none
module m;
endmodule
