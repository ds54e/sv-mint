`default_nettype none
module m;
endmodule
`default_nettype wire
