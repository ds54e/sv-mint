task t (
  inout logic a,
  input logic b,
  output logic c,
  ref logic d
);
endtask
