module parameter_violation #(
  parameter foo_value = 1,
  parameter BarValue = 2
) (); endmodule
