module header_missing;
endmodule
