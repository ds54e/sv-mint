`default_nettype none

module good;
endmodule

`default_nettype wire
