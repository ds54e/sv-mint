task t;
endtask
