module m;
  wire MyNet;
  wire MY_NET;
endmodule

