typedef enum int unsigned {
  off,
  on
} state_e;
