function logic f (logic a);
  return a;
endfunction
