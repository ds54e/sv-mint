`define GLOBAL_HELPER(x) (x)
