package FooPkg;
`define MACRO 1
endpackage : BarPkg

package AnotherPkg;
endpackage
