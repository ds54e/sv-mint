function logic f (input logic a);
  return 1'b0;
endfunction

