`default_nettype none

module port_names_lower_snake_violation(
  input logic Clk_i,
  output logic Data_o
);
endmodule

`default_nettype wire
