// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module net_lower_snake_violation;
  wire BadName;
endmodule

`default_nettype wire
