`define TEMP_MACRO(x) (x)
module macro_violation;
endmodule
