// SPDX-License-Identifier: Apache-2.0
// blank spacer

`timescale 1ns/1ps

module default_nettype_late;
  logic dummy0;
  logic dummy1;
  logic dummy2;
  logic dummy3;
  logic dummy4;
  logic dummy5;
  logic dummy6;
  logic dummy7;
  logic dummy8;
  logic dummy9;
  logic dummy10;
  logic dummy11;
  logic dummy12;
  logic dummy13;
  logic dummy14;
  logic dummy15;
  logic dummy16;
  logic dummy17;
  logic dummy18;
  logic dummy19;
  logic dummy20;
  logic dummy21;
endmodule

`default_nettype none

// forgot to reset to wire
