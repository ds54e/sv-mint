module my_module;
  `define MY_MODULE_MACRO
endmodule

