`default_nettype none

package pkg_with_define;
`define FOO 1
endpackage

`default_nettype wire
