module include_child;
  logic unused_signal;
endmodule
