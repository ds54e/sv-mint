module m;
  logic MyVar;
  logic MY_VAR;
endmodule

