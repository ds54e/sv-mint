module my_module;
  `define MACRO
endmodule

