`define UNUSED_MACRO 1

module macro_unused;
endmodule
