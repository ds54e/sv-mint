typedef logic [3:0] my_type_t;
