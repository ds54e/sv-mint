module m;
  logic a;
  always_comb begin
    a = 1'b1;
  end
endmodule
