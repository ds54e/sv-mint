module whitespace_violations;
	logic foo;
assign foo = 1'b0;  
endmodule
