// SPDX-License-Identifier: Apache-2.0
// Decl unused var compliant
`default_nettype none

module unused_var_compliant;

logic debug_shadow; // unused

endmodule

`default_nettype wire
