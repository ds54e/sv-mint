`default_nettype none

module module_name_matches_filename_good;
endmodule

`default_nettype wire
