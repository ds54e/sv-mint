module MyModule;
endmodule

module MY_MODULE;
endmodule
