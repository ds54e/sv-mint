task t (
  input a,
  output b
);
endtask
