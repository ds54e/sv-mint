automatic task t1;
endtask

static task t2;
endtask
