`default_nettype none

package pkg_one;
endpackage

package pkg_two;
endpackage

`default_nettype wire
