function acc_fn(input a_i, input b_i);
  acc_fn = a_i + b_i;
endfunction
