`default_nettype none
`define UNUSED_MACRO 1

module macro_unused;
endmodule

`default_nettype wire
