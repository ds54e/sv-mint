// Decl unused net violation
`default_nettype none

module unused_net_violation;

wire debug_tap;

endmodule

`default_nettype wire
