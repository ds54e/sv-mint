module m (
  input logic a,
  input logic b1, // reserved
  input logic b2, // used
  output logic c
);
  assign c = a;
endmodule

