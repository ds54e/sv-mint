module m #(
  parameter int my_param = 1,
  parameter int MY_PARAM = 1
);
endmodule
