`default_nettype none

module default_nettype_begins_with_none_good;
endmodule

`default_nettype wire
