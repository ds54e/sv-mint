module m #(
  localparam int MyParam = 1,
  localparam int MY_CONST = 1
);
endmodule
