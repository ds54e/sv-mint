﻿// SPDX-License-Identifier: Apache-2.0
module bom_crlf;
  wire [127:0] data_line_is_way_too_long_because_it_has_many_characters_which_should_break_rules_for_real_this_time;
endmodule
