`define MY_MACRO(a) a
