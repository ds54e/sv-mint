module not_bad;
endmodule
