// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module parameter_case_violation;
  parameter int data_width = 32;
endmodule

`default_nettype wire
