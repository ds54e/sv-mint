function automatic logic f1 (input logic a);
  return 1'b0;
endfunction

function static logic f2 (input logic a);
  return 1'b0;
endfunction

