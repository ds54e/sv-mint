function automatic f (input logic a);
  return 1'b0;
endfunction

