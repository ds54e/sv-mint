module m (
  inout logic my_port_1,
  input logic my_port_2,
  output logic my_port_3
);
endmodule
