`default_nettype none

typedef enum logic [1:0] {
  GOOD_ENUM_A,
  GOOD_ENUM_B
} good_enum_e;

module enum_type_names_lower_snake_e_good;
endmodule

`default_nettype wire
