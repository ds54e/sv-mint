`default_nettype none

package no_define_inside_package_good;
endpackage

`default_nettype wire
