module m;
  logic my_var;
  logic my_var$abc;
endmodule

