`include "include_child.sv"
module include_top;
endmodule
