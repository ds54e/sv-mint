// Decl unused net compliant
`default_nettype none

module unused_net_compliant;

wire debug_tap; // unused

endmodule

`default_nettype wire
