`default_nettype none

`define TEMP_MACRO(x) (x)
module macros_close_with_undef_bad;
endmodule

`default_nettype wire
