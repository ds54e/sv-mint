module m (
  inout logic a_io
  input logic b_i,
  output logic c_o
);
endmodule
