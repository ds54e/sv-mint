`default_nettype none

module net_lower_snake_ok;
  wire good_name;
  wire dollar_name;
endmodule

`default_nettype wire
