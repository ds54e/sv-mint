// Decl unused var violation
`default_nettype none

module unused_var_violation;

logic debug_shadow;

endmodule

`default_nettype wire
