module default_nettype_missing;
  logic a;
endmodule
