`default_nettype none

function automatic logic fn (
  input logic [1:0] a
);
  return 1'b0;
endfunction

`default_nettype wire
