program automatic main_program;
  initial begin
    $display("program block");
  end
endprogram
