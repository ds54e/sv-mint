module m #(
  parameter MyParam1 = 1,
  parameter MyParam2 = 1.0
);
endmodule
