`default_nettype none

module one_module_per_file_good;
endmodule

`default_nettype wire
