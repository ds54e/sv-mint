module m (
  inout logic a,
  input logic b,
  output logic c
);
endmodule

