`default_nettype none

module multiple_modules_ok;
endmodule

`default_nettype wire
