module m1 (
  inout logic MyPort1,
  input logic MyPort2,
  output logic MyPort3
);
endmodule

module m2 (
  inout logic MY_PORT_1,
  input logic MY_PORT_2,
  output logic MY_PORT_3
);
endmodule
