// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module module_filename_match_ok;
endmodule

`default_nettype wire
