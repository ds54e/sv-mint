`default_nettype none

`include "include_child.sv"
module include_top;
endmodule

`default_nettype wire
