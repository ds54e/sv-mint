function logic add(
  input logic a,
  input logic b
);
  return 1'b0;
endfunction
