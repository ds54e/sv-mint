task t (
  input logic a,
  output logic b
);
endtask
