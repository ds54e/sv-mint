`define MY_MACRO
