`default_nettype none

module foo;
endmodule

module bar;
endmodule

`default_nettype wire
