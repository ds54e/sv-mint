function logic add(
  input a,
  input b
);
  return 1'b0;
endfunction
