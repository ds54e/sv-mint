module foo_bar;
  `define FOO_BAR_LOCAL_MACRO(x) (x)
endmodule
