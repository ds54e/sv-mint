// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module single;
endmodule

`default_nettype wire
