`default_nettype none

typedef logic [3:0] good_type_t;

module typedef_names_lower_snake_t_good;
endmodule

`default_nettype wire
