`default_nettype none

module include_child;
  logic unused_signal;
endmodule

`default_nettype wire
