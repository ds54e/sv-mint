// SPDX-License-Identifier: Apache-2.0
// Decl unused param violation
`default_nettype none

module unused_param_violation #(
  parameter int EnableDbg = 0
) ();

endmodule

`default_nettype wire
