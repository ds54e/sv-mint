`default_nettype none

module module_filename_match_ok;
endmodule

`default_nettype wire
