`default_nettype none

module parameter_missing_type;
  parameter WIDTH = 4;
endmodule

`default_nettype wire
