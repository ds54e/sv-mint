module port_suffix_violation (
  input  logic clk,
  input  logic rst_n,
  output logic ready
);

endmodule
