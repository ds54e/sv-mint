`default_nettype none

`define badMacro 1

module macro_define_upper_violation;
endmodule

`default_nettype wire
