module m;
  wire a;
endmodule
