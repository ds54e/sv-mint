module m #(
  localparam MyParam1 = 1,
  localparam MyParam2 = 1.0
);
endmodule

