module m;
endmodule
