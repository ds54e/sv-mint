`default_nettype none

module wrong_name;
endmodule

`default_nettype wire
