// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module wrong_name;
endmodule

`default_nettype wire
