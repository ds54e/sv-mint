`default_nettype none

`define GOOD_MACRO 1

module macro_define_upper_ok;
endmodule

`default_nettype wire

`undef GOOD_MACRO
