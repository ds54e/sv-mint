module indent_violation;
   logic a;
   logic b;
`ifdef FOO
  logic c;
`endif
endmodule
