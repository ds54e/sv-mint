typedef logic [3:0] MyType_t;
typedef logic [3:0] MY_TYPE;
