`default_nettype none

module BadModuleName;
endmodule

`default_nettype wire
