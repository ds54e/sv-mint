function logic add(
  input logic a,
  b // missing direction
);
  return a + b;
endfunction
