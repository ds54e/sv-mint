`default_nettype none

package one_package_per_file_good;
endpackage

`default_nettype wire
