task t (
  logic a,
  logic b,
  logic c,
  logic d
);
endtask
