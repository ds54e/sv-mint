`default_nettype none

module port_names_suffix_violation(
  input logic clk,
  output logic data
);
endmodule

`default_nettype wire
