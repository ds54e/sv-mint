// SPDX-License-Identifier: Apache-2.0
`default_nettype none

module parameter_case_ok;
  parameter int DataWidth = 32;
  parameter int DATA_WIDTH = 16;
endmodule

`default_nettype wire
