`define my_macro
`define MyMacro
