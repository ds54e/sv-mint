`default_nettype none

typedef enum logic [1:0] {
  GoodValue,
  GOOD_VALUE
} enum_values_uppercase_good_e;

module enum_values_uppercase_good;
endmodule

`default_nettype wire
