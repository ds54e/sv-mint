`default_nettype none

module foo;
`define BAR 1
endmodule

`default_nettype wire
