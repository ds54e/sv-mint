class randomize_violation;
  function void run();
    req.randomize();
  endfunction
endclass
