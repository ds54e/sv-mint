module foo_bar;
  `define LOCAL_MACRO(x) (x)
endmodule
