`default_nettype wire

module default_nettype_wire;
endmodule
