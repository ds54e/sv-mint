module m # (
  parameter int MyParam = 1
);
endmodule
