`default_nettype none

module default_nettype_no_reset_violation;
endmodule
