module m #(
  localparam int my_const = 1
);
endmodule

