module m;
  wire my_net;
  wire my_net$abc;
endmodule
