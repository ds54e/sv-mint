typedef enum int unsigned {
  OFF,
  ON
} state_e;
