package function_scope_pkg;
function void helper();
endfunction
endpackage
