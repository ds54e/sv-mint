function logic f (input logic a);
  return a;
endfunction
