`default_nettype none

module parameter_range_only_violation;
  parameter [7:0] WIDTH = 8;
endmodule

`default_nettype wire
