module m #(
  localparam int unsigned MyParam1 = 1,
  localparam real MyParam2 = 1.0
);
endmodule

