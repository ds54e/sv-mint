module m (
  input logic a,
  output logic b
);
  assign b = 1'b1;
endmodule

