typedef enum int unsigned {
  OFF,
  ON
} state_1_e;

typedef enum int unsigned {
  Off,
  On
} state_2_e;
