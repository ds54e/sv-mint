`define DV_LOCAL_MACRO(x) (x)

module local_dv_macro;
endmodule

`undef DV_LOCAL_MACRO
