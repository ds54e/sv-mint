`default_nettype none

module disable_targets_fork_only_good;
endmodule

`default_nettype wire
