module sample(input logic clk);
  logic unused_var;
  logic net_unused;
  logic used_var;
  assign used_var = clk;
endmodule
