`define MY_MACRO(a) a
`undef MY_MACRO
