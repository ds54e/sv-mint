`default_nettype none

module default_nettype_ends_with_wire_good;
endmodule

`default_nettype wire
